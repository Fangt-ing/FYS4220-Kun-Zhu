library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity upCounter is
    port(
        sw
    );

end upCounter;

architecture upCount of upCounter is
    signal

    begin

end upCount;