library ieee;
context ieee.ieee_std_context;
use ieee.math_real.all;


entity system_top is
    port (
        clk   : in std_logic;
        arst_n : in std_logic;
        
    );
end entity;