library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;


package uart_rx_pakage is
    
end package;

package body uart_rx_pakage is
    
end package body;