component nios2_system is
    port (
    clk_clk       : in std_logic := 'X'; -- clk
    reset_reset_n : in std_logic := 'X'  -- reset_n

end component nios2_system;

u0 : component nios2_system
    port map(
        clk_clk       => CONNECTED_TO_clk_clk,      --   clk.clk
        reset_reset_n => CONNECTED_TO_reset_reset_n -- reset.reset_n
    )