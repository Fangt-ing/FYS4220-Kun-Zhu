��l i b r a r y   I E E E ;  
 u s e   I E E E . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
  
 e n t i t y   l a b 1   i s  
     p o r t   (  
             s w   :   i n   s t d _ l o g i c _ v e c t o r ( 9   d o w n t o   0 ) ;   - -   s l i d e   s w i t c h   a s   t h e   i n p u t s .  
             l e d   :   o u t   s t d _ l o g i c _ v e c t o r ( 9   d o w n t o   0 )   - -   l e d   a s   t h e   o u t p u t s .  
             ) ;  
         e n d   e n t i t y   l a b 1 ;  
  
 a r c h i t e c t u r e   t o p _ l e v e l   o f   l a b 1   i s  
  
 b e g i n  
         l e d   < =   s w ;  
 e n d   a r c h i t e c t u r e   t o p _ l e v e l ; 